module dff_reg(
    
    );