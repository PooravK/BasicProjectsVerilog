module register4bit(
    
    );