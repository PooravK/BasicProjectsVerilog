module basics;
  initial begin
    $display("Hello world");
    $finish;
  end
endmodule