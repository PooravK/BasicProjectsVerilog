module NotGate(input in, output out);
    assign out = !(in);
endmodule